module passthrough(input in,
                   output out);

   assign out = in;

endmodule
